library verilog;
use verilog.vl_types.all;
entity key_to_seg7_vlg_vec_tst is
end key_to_seg7_vlg_vec_tst;
